module JumpControl (
	input				[4:0]		opcode_i
);

endmodule	